module tb;
    reg [0:1] Select;
    reg [0:3] AccountNumber;
    reg [0:9] Balance;
    wire [0:9] Output;
endmodule